* Minimum Output Voltage for proper working of Current Mirror

VDD 3 0 DC 5v
VDS 2 0 DC 5v
M1 1 1 0 0 NMOS12 W=5u L=1u
M2 2 1 0 0 NMOS12 W=5u L=1u
IREF 3 1 20u
.MODEL NMOS12 NMOS(kp=200u LAMBDA=0.01 VTO=0.4)
.DC VDS 0 1 0.01
.op
.PROBE
.END



