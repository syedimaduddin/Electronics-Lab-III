* Simulation of Common Emitter Amplifier

Vin 1 0 sin(0 10m 1k)
C1 1 2 10uF
Rb 2 3 10k
R1 4 2 12k
R2 2 0 1k
Vcc 4 0 DC 15v
Rc 4 5 1k
Q1 5 3 0 Q2N2222
.model Q2N2222	NPN(Is=14.34f Xti=3 Eg=1.11 Vaf=74.03 Bf=255.9 Ne=1.307
+		Ise=14.34f Ikf=.2847 Xtb=1.5 Br=6.092 Nc=2 Isc=0 Ikr=0 Rc=1
+		Cjc=7.306p Mjc=.3416 Vjc=.75 Fc=.5 Cje=22.01p Mje=.377 Vje=.75
+		Tr=46.91n Tf=411.1p Itf=.6 Vtf=1.7 Xtf=3 Rb=10)
*		National	pid=19		case=TO18
*		88-09-07 bam	creation
.TRAN 0.1u 5m
.PROBE
.END

