
*----------------------------------------
* Syed Imaduddin_20ELB124
*----------------------------------------

Vin 1 0 sin(0 5v 10KHz)
C1 1 2 10uF
D1 0 2 DIN914
R1 2 0 1k
.MODEL DIN914 D()
.TRAN 0.1MS 0.5MS 
.PROBE
.END
*----------------------------------------



