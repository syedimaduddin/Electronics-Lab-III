
*----------------------------------------
* Syed Imaduddin_20ELB124
*----------------------------------------

* Diode Characteristics

Vin 1 0 2v
R1 1 2 550
D1 2 0 D1N914
.MODEL D1N914 D()
.DC lin Vin 0 2v 0.1v
.PROBE
.END

*----------------------------------------
