
*----------------------------------------
* Syed Imaduddin_20ELB124
*----------------------------------------

Vin 1 0 sin(0 5v 5KHz)
R1 1 2 1k
DA 2 3 DIN914
.MODEL DIN914 D()
V1 3 0 2v
.TRAN 0.1MS 1MS
.PROBE
.END

*----------------------------------------


