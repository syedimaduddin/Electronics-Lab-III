* MOS Current Mirror for Different current ratios

VDD 3 0 DC 5v
RL 3 2 1k
M1 1 1 0 0 NMOS12 W=5u L=1u
M2 2 1 0 0 NMOS12 W={W2} L=1u
IREF 3 1 20u
.MODEL NMOS12 NMOS(kp=200u LAMBDA=0 VTO=0.5)
.PARAM W2=1
.STEP PARAM W2 LIST 5u 10u 20u
.DC IREF 0 50u 1u 
.PROBE
.END


