
*----------------------------------------
* Syed Imaduddin_20ELB124
*----------------------------------------

Vin 1 0 sin(0 10v 10KHz)
R1 1 2 1k
D1 2 3 DIN914
V1 3 0 5v
D2 4 2 DIN914
V2 0 4 5v
.MODEL DIN914 D()
.TRAN 0.1MS 0.5MS
.PROBE
.END
*----------------------------------------


